`include "design.v"
`include "add.sv"
`include "addG.sv"
`include "sub.sv"
`include "subG.sv"
`include "mul.sv"
`include "div.sv"
`include "comparator.sv"
`include "div_fsmLS.sv"
`include "mux16to1.sv"
`include "mux4to1.sv"
`include "demux1to16.sv"
